library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity image is
    port(
      --  clk: in std_logic;
        addr: in unsigned(4 downto 0);
        data: out std_logic_vector(0 to 127)

    );
end image;

architecture content of image is
    type rom_type is array(0 to 31) of std_logic_vector(127 downto 0);
    constant IMG: rom_type :=
    (
        "00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000111100000000000000000000000000000000001111000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000111000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000110000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000",
        "00000000000000000000000000011000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000",
        "00000000000000000000000000100000000000000111111111000000000000111111111000000000000001000000000000000000000000000000000000000000",
        "00000000000000000000000001000000000111110000000000111000000111000000000011111000000000100000000000000000000000000000000000000000",
        "00000000000000000000000010000000110000000000000000000110011000000000000000000011000000010000000000000000000000000000000000000000",
		  "00000000000011111110000100000001000000000000000000000000000000000000000000000000100000001000011111110000000000000000000000000000",
        "00000000001000000001100100000010000111111111110000000000000000000011111111111000010000001001100000000100000000000000000000000000",
        "00000000010000000000110100000100000000000000000000000000000000000000000000000000001000001011000000000010000000000000000000000000",
        "00000000010000000000011100001000000000000000000000000000000000000000000000000000000100001110000000000010000000000000000000000000",
        "00000000010000000000000100010000000000000000000000000000000000000000000000000000000010001000000000000010000000000000000000000000",
        "00000000010000000000000100010000000000000111100000000000000000000001111000000000000010001000000000000010000000000000000000000000",
        "00000000010000000000000100010000000000000111100000000000000000000001111000000000000010001000000000000010000000000000000000000000",
        "00000000010000000000000100010000000000000000000000000000000000000000000000000000000010001000000000000010000000000000000000000000",
		  "00000000010000000000001100010000000000000000000000000000000000000000000000000000000010001100000000000010000000000000000000000000",
        "00000000001000000001100100010000000000000000000000000000000000000000000000000000000010001001100000000100000000000000000000000000",
        "00000000000011111110000100010000000000000001111000000111111000001111100000000000000010001000011111110000000000000000000000000000",
        "00000000000000000000000100011000000000000010000000000011110000000000010000010000000110001000000000000000000000000000000000000000",
        "00000000000000000000000100000111000000000100000000000000000000000000001010000000111000001000000000000000000000000000000000000000",
        "00000000000000000000000100000000111100000100000000000000000000000000001000001111000000001000000000000000000000000000000000000000",
        "00000000000000000000000001100000000011111100000000000000000000000000001111110000000001100000000000000000000000000000000000000000",
        "00000000000000000000000000011000000000000100000000000000000000000000001000000000000110000000000000000000000000000000000000000000",
		  "00000000000000000000000000000110000000000100000000000000000000000000001000000000011000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000111000000100000000000000000000000000001000000111000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000111000100000000000000000000000000001000111000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000011101000000000000000000000000101110000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000010100000000000000000000001010000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000101111111111111111111101000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000"
		  
     );
begin
     data <= IMG(to_integer(addr));
end content;

