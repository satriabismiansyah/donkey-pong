library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity bar_rom is
    port(
        clk: in std_logic;
        addr: in unsigned(2 downto 0);
        data: out std_logic_vector(0 to 127); 
		  
		  addr2: in unsigned(2 downto 0);
        data2: out std_logic_vector(0 to 127)
    );
end bar_rom;

architecture content of bar_rom is
    type rom_type is array(0 to 7) of std_logic_vector(127 downto 0);
    constant BAR: rom_type :=
    (
        "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
        "11000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011",
        "11000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011",
        "11000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011",
        "11000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011",
        "11000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011",
        "11000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011",
        "11000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011"
    );
    signal addr_reg: unsigned(2 downto 0);
    signal addr_reg2: unsigned(2 downto 0);
begin
    process(clk)
    begin
        if rising_edge(clk) then
            addr_reg <= addr;
        end if;
    end process;      
	 
	  process(clk)
    begin
        if rising_edge(clk) then
            addr_reg2 <= addr2;
        end if;
    end process;            
    data <= BAR(to_integer(addr_reg));
    data2 <= BAR(to_integer(addr_reg2));
end content;

